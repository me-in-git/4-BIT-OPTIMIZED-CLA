// Pragnya_2023102067 
module xor_sum (
    output xor_z,
    input cin, k
);
    assign xor_z = cin ^ k;  // XOR for sum computation
endmodule
