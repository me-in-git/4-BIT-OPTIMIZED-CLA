* SPICE3 file created from xor.ext - technology: scmos

.option scale=1u

M1000 inv_0/op a vdd inv_0/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=360 ps=184
M1001 inv_0/op a gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=121 ps=79
M1002 inv_1/op b vdd inv_1/w_0_6# pfet w=12 l=2
+  ad=60 pd=34 as=0 ps=0
M1003 inv_1/op b gnd Gnd nfet w=6 l=2
+  ad=30 pd=22 as=0 ps=0
M1004 op inv_0/op a_10_10# w_n3_4# pfet w=24 l=2
+  ad=192 pd=64 as=432 ps=180
M1005 vdd a_18_0# a_10_10# w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 gnd inv_1/op a_38_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=96 ps=40
M1007 a_10_10# inv_1/op op w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_10_n43# a_8_n46# gnd Gnd nfet w=12 l=2
+  ad=96 pd=40 as=0 ps=0
M1009 a_38_n43# inv_0/op op Gnd nfet w=12 l=2
+  ad=0 pd=0 as=120 ps=68
M1010 op a_18_n46# a_10_n43# Gnd nfet w=12 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_10_10# a_8_1# vdd w_n3_4# pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
C0 inv_1/op a_8_n46# 0.18fF
C1 w_n3_4# a_8_1# 2.62fF
C2 inv_1/op b 0.20fF
C3 inv_1/op inv_0/op 0.18fF
C4 vdd inv_0/w_0_6# 0.85fF
C5 inv_1/w_0_6# vdd 0.85fF
C6 b a_8_n46# 0.11fF
C7 inv_0/op w_n3_4# 2.62fF
C8 w_n3_4# a_18_0# 2.62fF
C9 inv_0/op a_8_n46# 0.18fF
C10 inv_0/op a 0.61fF
C11 inv_0/op b 0.41fF
C12 inv_1/w_0_6# inv_1/op 0.85fF
C13 a_10_10# w_n3_4# 4.37fF
C14 inv_1/op op 0.36fF
C15 inv_1/op a_18_n46# 0.18fF
C16 a_10_10# a_18_0# 0.18fF
C17 a inv_0/w_0_6# 2.62fF
C18 w_n3_4# op 0.85fF
C19 inv_1/w_0_6# b 3.61fF
C20 inv_0/op inv_0/w_0_6# 0.85fF
C21 vdd w_n3_4# 1.69fF
C22 vdd b 0.47fF
C23 inv_0/op op 0.18fF
C24 inv_0/op a_18_n46# 0.18fF
C25 gnd a 0.47fF
C26 inv_1/op w_n3_4# 2.62fF
C27 a_18_n46# Gnd 7.54fF
C28 a_8_n46# Gnd 7.78fF
C29 op Gnd 0.99fF
C30 a_18_0# Gnd 1.11fF
C31 a_8_1# Gnd 0.87fF
C32 inv_1/op Gnd 21.28fF
C33 b Gnd 12.44fF
C34 gnd Gnd 12.88fF
C35 inv_0/op Gnd 21.14fF
C36 vdd Gnd 8.04fF
C37 a Gnd 11.02fF
